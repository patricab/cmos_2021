.include ../models/ptm_130.spi
.include ../lib/SUN_TRIO_GF130N.spi

.include comp.cir

.option TNOM=27 GMIN=1e-20

* Main circuit
.subckt pixel_sensor VBN1 RAMP RESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

*** Subcircuit calls
* XS1 VRESET VSTORE ERASE EXPOSE VDD VSS SENSOR
* XC1 VCMP_OUT VSTORE VRAMP VDD VSS COMP
XCM VDD VSS PG RAMP VBN1 DATA
* XM1 READ VCMP_OUT DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS MEMORY
.ends
