.include ../models/ptm_130_ngspice.spi
.include ../lib/SUN_TR_GF130N.spi
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6

* Analog parameters
* .param VDD = 1.5

* Sources
VDD VDD VSS dc 1.5
VSS VSS 0 dc 0
VPG VPG 0 dc 1
VRAMP VRAMP 0 dc 0

* Bias
IPB1 0 VBN1 dc 1u
XMNB0 VBN1 VBN1 VSS VSS NCHCM2

* DUT
.include pixelSensor.cir
XDUT VDD VSS VPG VRAMP VBN1 VOUT COMP
* .subckt COMP VDD VSS PG RAMP VBN1 OUT

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
* Sweeps
* dc VPG 0 2 0.001
dc VRAMP 0 2 0.001

* Plot/write to file
* plot V(VOUT) V(VPG) V(VRAMP)
plot V(VOUT) 
* hardcopy plot.ps V(VOUT)
.endc
.end