.include ../models/ptm_130.spi
.include ../lib/SUN_TRIO_GF130N.spi

* Comparator 
.subckt COMP VPG VRAMP OUT VBN1 VDD VSS 
VBT VBT 0 dc 0.3

* PMOS Current Mirror
MP1 VCM VCM VDD VDD pmos w=0.5u l=0.5u
MP2 CMP VCM VDD VDD pmos w=0.5u l=0.5u

* Differential amplifier
MN1 VCM VPG VB VSS nmos w=0.5u l=0.5u 
MN2 CMP VRAMP VB VSS nmos w=0.5u l=0.5u

* Bias transistor
XB1 VB VBN1 VSS VSS NCHCM2

* Common source amplifier
MP3 VDD CMP VINV VSS pmos l=0.5u w=0.5u
MN4 VINV VBT VSS VSS nmos l=0.5u w=0.5u

* Inverter
MP4 VDD VINV OUT VDD pmos L=0.5u W=0.5u 
MN5 OUT VINV VSS VSS nmos L=0.5u W=0.5u

* Output capacitor
CL OUT VSS 1p
.ends
