.include ../models/ptm_130.spi
.include ../lib/SUN_TRIO_GF130N.spi

.include comp.cir
.include sens.cir

.option TNOM=27 GMIN=1e-20

* Main circuit
.subckt pixel_sensor VBN1 VRAMP VRESET ERASE EXPOSE READ
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

*** Subcircuit calls
* Sensor
XSENS VRESET PG ERASE EXPOSE VDD VSS sens
* .subckt sens VRESET VSTORE ERASE EXPOSE VDD VSS

* Comparator
XCMP PG VRAMP VBN1 CMP VDD VSS COMP
* .subckt COMP PG RAMP VBN1 OUT VDD VSS

* Memory
XMEM READ CMP DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS 
+ MEMORY
.ends

* Copied from dicex
.SUBCKT MEMORY READ VCMP_OUT
+ DATA_7 DATA_6 DATA_5 DATA_4 DATA_3 DATA_2 DATA_1 DATA_0 VDD VSS

XM1 VCMP_OUT DATA_0 READ VSS MEMCELL
XM2 VCMP_OUT DATA_1 READ VSS MEMCELL
XM3 VCMP_OUT DATA_2 READ VSS MEMCELL
XM4 VCMP_OUT DATA_3 READ VSS MEMCELL
XM5 VCMP_OUT DATA_4 READ VSS MEMCELL
XM6 VCMP_OUT DATA_5 READ VSS MEMCELL
XM7 VCMP_OUT DATA_6 READ VSS MEMCELL
XM8 VCMP_OUT DATA_7 READ VSS MEMCELL
.ENDS

.SUBCKT MEMCELL CMP DATA READ VSS
M1 VG CMP DATA VSS nmos  w=0.2u  l=0.13u
M2 DATA READ DMEM VSS nmos  w=0.4u  l=0.13u
M3 DMEM VG VSS VSS nmos  w=1u  l=0.13u
C1 VG VSS 1p
.ENDS